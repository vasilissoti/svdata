module TestModule
( output var signed [FOO-1:0] a, b
, output var logic signed c, reg signed d
, output logic signed e [DOO-1:0]
, output integer signed f
);
endmodule