module Boo
( input tri a
, input reg b
, output signed c, d
, output logic signed e
);
endmodule
