module mh20(ref x [5:0], y);
endmodule