module Koo
( [5:0] x
);
endmodule
