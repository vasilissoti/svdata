module mh4 (input x);
endmodule