module TestModule
( output [FOO-1:0] a, b
, output wire logic [FOO-1:0] c, wire reg d
, output wire string e
, output tri integer unsigned f
);
endmodule