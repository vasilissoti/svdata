module mh19(ref [5:0] x, y);
endmodule