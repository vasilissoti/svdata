module mh18(output signed [5:0] x, integer y);
endmodule