package TestPackage;
  /*pre*/ parameter /*kw/ty*/ a /*post*/ = /*eq/val*/ 1 /* post */;
  /*pre*/ parameter /*kw/ty*/ b /* id/eq */ = /*eq/val*/ 5 /* post */;
  /*pre*/ parameter /*kw/ty*/ int /*ty/id*/ c /*post*/ = /*eq/val*/ 3 /* post */;
  /*pre*/ parameter /*kw/ty*/ int /*ty/id*/ d /*id/eq*/ = /*eq/val*/ 2 /*post*/;
  /*pre*/ localparam /*kw/ty*/ e /* id/eq */ = /*eq/val*/ 5 /* post */;
  /*pre*/ localparam /*kw/ty*/ int /*ty/id*/ f /*id/eq*/ = /*eq/val*/ 5 /*post*/;
endpackage