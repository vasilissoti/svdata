module mh8 (output var x);
endmodule