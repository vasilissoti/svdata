module TestModule
( output var signed [FOO-1:0] a [FOO] [FOO-1:0], b
, output var logic signed c, reg signed d
, output logic signed e [FOO-1:0]
, output integer signed f
);
endmodule