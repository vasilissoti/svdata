module M #() ();
  I #(.A(A)) u_I [B-1:0] (.a());
endmodule
