module TestModule
( output tri my_enum_t d
, output wire my_struct_t e, f
);
endmodule