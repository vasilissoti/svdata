module TestModule
( output var [FOO-1:0] a [FOO] [FOO-1:0], b
, output var logic c, reg d
, output logic unsigned e [FOO-1:0]
, output string f
, output integer unsigned g
);
endmodule