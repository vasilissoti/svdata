module mh6 (input var integer x);
endmodule