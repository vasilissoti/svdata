module TestModule
#(parameter signed a = 8'b10101010, 
  parameter logic signed [3:0] b = 4'b1000, c [4:0],
  parameter my_struct d,
  parameter e = 7.5, f = 5)
(); 
endmodule