module TestModule
( input [FOO-1:0] a, b
, input wire [FOO-1:0] c [FOO] [FOO-1:0], reg d
, input logic e [FOO-1:0]
, input string f
, input tri integer unsigned g
);
endmodule