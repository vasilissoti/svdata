module mh0 (wire x);
endmodule