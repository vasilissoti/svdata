module mh15([5:0] x, wire y);
endmodule