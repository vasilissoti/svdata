module testmodule(
    input a, b,
    output a2, b2
  );

  bar test0 (.a(a2[i]), .b(b2[k])); 
  bar test1 (.a(a2[i]), .b(b2[k])); 

endmodule
