module TestModule
( input var my_enum_t d
, input var my_struct_t e, f
);
endmodule