module TestModule
#(integer signed a = 8'b10101010, 
  logic signed [3:0] b = 4'b1000, c [4:0],
  real e = 7.5, 
  integer f = 5)
(); 
endmodule