module mh13(wire x, y[7:0]);
endmodule