module mh14(integer x, signed [5:0] y);
endmodule