module mh10(output integer x);
endmodule