module mh11(ref [5:0] x);
endmodule