module TestModule
( output var [FOO-1:0] a, b
, output var logic c, reg d
, output logic unsigned e [DOO-1:0]
, output string f
, output integer unsigned g
);
endmodule