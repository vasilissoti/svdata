module mh5 (input var x);
endmodule