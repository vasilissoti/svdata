module TestModule
( input my_enum_t d
, input wire my_struct_t e, f
);
endmodule