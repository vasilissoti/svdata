module Doo
( input var string tmp
, input int signed a, logic b
, output wire signed c, unsigned d
);
endmodule
