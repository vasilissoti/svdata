module TestModule
#(localparam signed a = 8'b10101010, 
  localparam logic signed [3:0] b = 4'b1000, c [4:0],
  localparam my_struct d,
  localparam e = 7.5, f = 5)
(); 
endmodule