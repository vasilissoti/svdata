package P_integralDataTypes; // {{{
  localparam shortint shortint_0 = 0;
  localparam shortint shortint_1 = 1;
  localparam shortint shortint_2 = -1;
  localparam shortint shortint_3 = 123;
  localparam shortint shortint_4 = 16'h5555;
  localparam shortint shortint_5 = 'h5556;
  localparam shortint shortint_6 = 'sh5557;
  localparam shortint shortint_7 = -16'h5558;
  localparam shortint shortint_8 = -'h5559;
  localparam shortint shortint_9 = -'sh5560;
  localparam shortint shortint_10 = 16'd5555;
  localparam shortint shortint_11 = 'd5556;
  localparam shortint shortint_12 = 'sd5557;
  localparam shortint shortint_13 = -16'd5558;
  localparam shortint shortint_14 = -'d5559;
  localparam shortint shortint_15 = -'sd5560;
  localparam shortint shortint_16 = '0;
  localparam shortint shortint_17 = '1;
  localparam shortint unsigned shortint_unsigned_0 = 0;
  localparam shortint unsigned shortint_unsigned_1 = 1;
  localparam shortint unsigned shortint_unsigned_2 = -1;
  localparam shortint unsigned shortint_unsigned_3 = 123;
  localparam shortint signed shortint_signed_0 = 0;
  localparam shortint signed shortint_signed_1 = 1;
  localparam shortint signed shortint_signed_2 = -1;
  localparam shortint signed shortint_signed_3 = 123;

  localparam int int_0 = 0;
  localparam int int_1 = 1;
  localparam int int_2 = -1;
  localparam int int_3 = 123;
  localparam int int_4 = 32'h5555_0505;
  localparam int int_5 = 'h5556;
  localparam int int_6 = 'sh5557;
  localparam int int_7 = -32'h5558_0505;
  localparam int int_8 = -'h5559;
  localparam int int_9 = -'sh5560;
  localparam int int_10 = 32'd5555;
  localparam int int_11 = 'd5556;
  localparam int int_12 = 'sd5557;
  localparam int int_13 = -32'd5558;
  localparam int int_14 = -'d5559;
  localparam int int_15 = -'sd5560;
  localparam int int_16 = '0;
  localparam int int_17 = '1;
  localparam int unsigned int_unsigned_0 = 0;
  localparam int unsigned int_unsigned_1 = 1;
  localparam int unsigned int_unsigned_2 = -1;
  localparam int unsigned int_unsigned_3 = 123;
  localparam int signed int_signed_0 = 0;
  localparam int signed int_signed_1 = 1;
  localparam int signed int_signed_2 = -1;
  localparam int signed int_signed_3 = 123;

  localparam longint longint_0 = 0;
  localparam longint longint_1 = 1;
  localparam longint longint_2 = -1;
  localparam longint longint_3 = 123;
  localparam longint longint_4 = 64'h5555_0505_0505_0505;
  localparam longint longint_5 = 'h5556;
  localparam longint longint_6 = 'sh5557;
  localparam longint longint_7 = -64'h5558_0505_0505_0505;
  localparam longint longint_8 = -'h5559;
  localparam longint longint_9 = -'sh5560;
  localparam longint longint_10 = 64'd5555;
  localparam longint longint_11 = 'd5556;
  localparam longint longint_12 = 'sd5557;
  localparam longint longint_13 = -64'd5558;
  localparam longint longint_14 = -'d5559;
  localparam longint longint_15 = -'sd5560;
  localparam longint longint_16 = '0;
  localparam longint longint_17 = '1;
  localparam longint unsigned longint_unsigned_0 = 0;
  localparam longint unsigned longint_unsigned_1 = 1;
  localparam longint unsigned longint_unsigned_2 = -1;
  localparam longint unsigned longint_unsigned_3 = 123;
  localparam longint signed longint_signed_0 = 0;
  localparam longint signed longint_signed_1 = 1;
  localparam longint signed longint_signed_2 = -1;
  localparam longint signed longint_signed_3 = 123;

  localparam byte byte_0 = 0;
  localparam byte byte_1 = 1;
  localparam byte byte_2 = -1;
  localparam byte byte_3 = 123;
  localparam byte byte_4 = 8'h55;
  localparam byte byte_5 = 'h56;
  localparam byte byte_6 = 'sh57;
  localparam byte byte_7 = -8'h58;
  localparam byte byte_8 = -'h59;
  localparam byte byte_9 = -'sh60;
  localparam byte byte_10 = 8'd55;
  localparam byte byte_11 = 'd56;
  localparam byte byte_12 = 'sd57;
  localparam byte byte_13 = -8'd58;
  localparam byte byte_14 = -'d59;
  localparam byte byte_15 = -'sd60;
  localparam byte byte_16 = '0;
  localparam byte byte_17 = '1;
  localparam byte unsigned byte_unsigned_0 = 0;
  localparam byte unsigned byte_unsigned_1 = 1;
  localparam byte unsigned byte_unsigned_2 = -1;
  localparam byte unsigned byte_unsigned_3 = 123;
  localparam byte signed byte_signed_0 = 0;
  localparam byte signed byte_signed_1 = 1;
  localparam byte signed byte_signed_2 = -1;
  localparam byte signed byte_signed_3 = 123;

  localparam bit bit_0 = 1'b0;
  localparam bit bit_1 = 1'b1;
  localparam bit bit_2 = '0;
  localparam bit bit_3 = '1;
  localparam bit unsigned bit_unsigned_0 = 1'b0;
  localparam bit unsigned bit_unsigned_1 = 1'b1;
  localparam bit signed bit_signed_0 = 1'b0;
  localparam bit signed bit_signed_1 = 1'b1;

  localparam logic logic_0 = 1'b0;
  localparam logic logic_1 = 1'b1;
  localparam logic logic_2 = '0;
  localparam logic logic_3 = '1;
  localparam logic logic_4 = 1'bX;
  localparam logic logic_5 = 1'bZ;
  localparam logic logic_6 = 'X;
  localparam logic logic_7 = 'Z;
  localparam logic logic_8 = -1;
  localparam logic logic_9 = 'sd57;
  localparam logic logic_10 = -8'd58;
  localparam logic logic_11 = -'sh60;
  localparam logic unsigned logic_unsigned_0 = 1'b0;
  localparam logic unsigned logic_unsigned_1 = 1'b1;
  localparam logic signed logic_signed_0 = 1'b0;
  localparam logic signed logic_signed_1 = 1'b1;

  localparam reg reg_0 = 1'b0;
  localparam reg reg_1 = 1'b1;
  localparam reg reg_2 = '0;
  localparam reg reg_3 = '1;
  localparam reg reg_4 = 1'bX;
  localparam reg reg_5 = 1'bZ;
  localparam reg reg_6 = 'X;
  localparam reg reg_7 = 'Z;
  localparam reg reg_8 = -1;
  localparam reg reg_9 = 'sd57;
  localparam reg reg_10 = -8'd58;
  localparam reg reg_11 = -'sh60;
  localparam reg unsigned reg_unsigned_0 = 1'b0;
  localparam reg unsigned reg_unsigned_1 = 1'b1;
  localparam reg signed reg_signed_0 = 1'b0;
  localparam reg signed reg_signed_1 = 1'b1;

  localparam integer integer_0 = 0;
  localparam integer integer_1 = 1;
  localparam integer integer_2 = -1;
  localparam integer integer_3 = 123;
  localparam integer integer_4 = 32'h5555_0505;
  localparam integer integer_5 = 'h5556;
  localparam integer integer_6 = 'sh5557;
  localparam integer integer_7 = -32'h5558_0505;
  localparam integer integer_8 = -'h5559;
  localparam integer integer_9 = -'sh5560;
  localparam integer integer_10 = 32'd5555;
  localparam integer integer_11 = 'd5556;
  localparam integer integer_12 = 'sd5557;
  localparam integer integer_13 = -32'd5558;
  localparam integer integer_14 = -'d5559;
  localparam integer integer_15 = -'sd5560;
  localparam integer integer_16 = '0;
  localparam integer integer_17 = '1;
  localparam integer integer_18 = 'X;
  localparam integer integer_19 = 'Z;
  localparam integer integer_20 = {8{4'b01XZ}};
  localparam integer unsigned integer_unsigned_0 = 0;
  localparam integer unsigned integer_unsigned_1 = 1;
  localparam integer unsigned integer_unsigned_2 = -1;
  localparam integer unsigned integer_unsigned_3 = 123;
  localparam integer signed integer_signed_0 = 0;
  localparam integer signed integer_signed_1 = 1;
  localparam integer signed integer_signed_2 = -1;
  localparam integer signed integer_signed_3 = 123;

  localparam time time_0 = 0;
  localparam time time_1 = 1;
  localparam time time_2 = -1;
  localparam time time_3 = 123;
  localparam time time_4 = 64'h5555_0505_0505_0505;
  localparam time time_5 = 'h5556;
  localparam time time_6 = 'sh5557;
  localparam time time_7 = -64'h5558_0505_0505_0505;
  localparam time time_8 = -'h5559;
  localparam time time_9 = -'sh5560;
  localparam time time_10 = 64'd5555;
  localparam time time_11 = 'd5556;
  localparam time time_12 = 'sd5557;
  localparam time time_13 = -64'd5558;
  localparam time time_14 = -'d5559;
  localparam time time_15 = -'sd5560;
  localparam time time_16 = '0;
  localparam time time_17 = '1;
  localparam time time_18 = 'X;
  localparam time time_19 = 'Z;
  localparam time time_20 = {16{4'b01XZ}};
  localparam time unsigned time_unsigned_0 = 0;
  localparam time unsigned time_unsigned_1 = 1;
  localparam time unsigned time_unsigned_2 = -1;
  localparam time unsigned time_unsigned_3 = 123;
endpackage // }}} P_integralDataTypes

package P_integralNonVectorUnpacked; // {{{
  localparam shortint shortint_0 [3] = '{1, 2, 3};
  localparam shortint shortint_1 [3] = '{-1, -2, -3};
  localparam shortint shortint_2 [3] = '{'1, '0, '1};
  localparam shortint unsigned shortint_unsigned_0 [3] = '{1, 2, 3};
  localparam shortint unsigned shortint_unsigned_1 [3] = '{-1, -2, -3};
  localparam shortint unsigned shortint_unsigned_2 [3] = '{'1, '0, '1};
  localparam shortint signed shortint_signed_0 [3] = '{1, 2, 3};
  localparam shortint signed shortint_signed_1 [3] = '{-1, -2, -3};
  localparam shortint signed shortint_signed_2 [3] = '{'1, '0, '1};

  localparam int int_0 [3] = '{1, 2, 3};
  localparam int int_1 [3] = '{-1, -2, -3};
  localparam int int_2 [3] = '{'1, '0, '1};
  localparam int unsigned int_unsigned_0 [3] = '{1, 2, 3};
  localparam int unsigned int_unsigned_1 [3] = '{-1, -2, -3};
  localparam int unsigned int_unsigned_2 [3] = '{'1, '0, '1};
  localparam int signed int_signed_0 [3] = '{1, 2, 3};
  localparam int signed int_signed_1 [3] = '{-1, -2, -3};
  localparam int signed int_signed_2 [3] = '{'1, '0, '1};

  localparam longint longint_0 [3] = '{1, 2, 3};
  localparam longint longint_1 [3] = '{-1, -2, -3};
  localparam longint longint_2 [3] = '{'1, '0, '1};
  localparam longint unsigned longint_unsigned_0 [3] = '{1, 2, 3};
  localparam longint unsigned longint_unsigned_1 [3] = '{-1, -2, -3};
  localparam longint unsigned longint_unsigned_2 [3] = '{'1, '0, '1};
  localparam longint signed longint_signed_0 [3] = '{1, 2, 3};
  localparam longint signed longint_signed_1 [3] = '{-1, -2, -3};
  localparam longint signed longint_signed_2 [3] = '{'1, '0, '1};

  localparam byte byte_0 [3] = '{1, 2, 3};
  localparam byte byte_1 [3] = '{-1, -2, -3};
  localparam byte byte_2 [3] = '{'1, '0, '1};
  localparam byte unsigned byte_unsigned_0 [3] = '{1, 2, 3};
  localparam byte unsigned byte_unsigned_1 [3] = '{-1, -2, -3};
  localparam byte unsigned byte_unsigned_2 [3] = '{'1, '0, '1};
  localparam byte signed byte_signed_0 [3] = '{1, 2, 3};
  localparam byte signed byte_signed_1 [3] = '{-1, -2, -3};
  localparam byte signed byte_signed_2 [3] = '{'1, '0, '1};

  localparam integer integer_0 [3] = '{1, 2, 3};
  localparam integer integer_1 [3] = '{-1, -2, -3};
  localparam integer integer_2 [3] = '{'1, '0, '1};
  localparam integer integer_3 [4] = '{'0, '1, 'X, 'Z};
  localparam integer unsigned integer_unsigned_0 [3] = '{1, 2, 3};
  localparam integer unsigned integer_unsigned_1 [3] = '{-1, -2, -3};
  localparam integer unsigned integer_unsigned_2 [3] = '{'1, '0, '1};
  localparam integer unsigned integer_unsigned_3 [4] = '{'0, '1, 'X, 'Z};
  localparam integer signed integer_signed_0 [3] = '{1, 2, 3};
  localparam integer signed integer_signed_1 [3] = '{-1, -2, -3};
  localparam integer signed integer_signed_2 [3] = '{'1, '0, '1};
  localparam integer signed integer_signed_3 [4] = '{'0, '1, 'X, 'Z};

  localparam time time_0 [3] = '{1, 2, 3};
  localparam time time_1 [3] = '{-1, -2, -3};
  localparam time time_2 [3] = '{'1, '0, '1};
  localparam time time_3 [4] = '{'0, '1, 'X, 'Z};
  localparam time unsigned time_unsigned_0 [3] = '{1, 2, 3};
  localparam time unsigned time_unsigned_1 [3] = '{-1, -2, -3};
  localparam time unsigned time_unsigned_2 [3] = '{'1, '0, '1};
  localparam time unsigned time_unsigned_3 [4] = '{'0, '1, 'X, 'Z};
  localparam time signed time_signed_0 [3] = '{1, 2, 3};
  localparam time signed time_signed_1 [3] = '{-1, -2, -3};
  localparam time signed time_signed_2 [3] = '{'1, '0, '1};
  localparam time signed time_signed_3 [4] = '{'0, '1, 'X, 'Z};
endpackage // }}} P_integralNonVectorUnpacked

package P_integralVectorPacked; // {{{
  localparam bit [3:0] bit_0 = 4'b0101;
  localparam bit [3:0] bit_1 = 4'd5;
  localparam bit [3:0] bit_2 = 5;
  localparam bit [3:0] bit_3 = '0;
  localparam bit [3:0] bit_4 = '1;
  localparam bit [2:0][3:0] bit_5 = '0;
  localparam bit [2:0][3:0] bit_6 = '1;
  localparam bit [2:0][3:0] bit_7 = '{1, 2, 3};
  localparam bit [2:0][3:0] bit_8 = {4'd1, 4'd2, 4'd3};
  localparam bit unsigned [3:0] bit_unsigned_0 = 4'b0101;
  localparam bit unsigned [3:0] bit_unsigned_1 = 4'd5;
  localparam bit unsigned [3:0] bit_unsigned_2 = 5;
  localparam bit unsigned [3:0] bit_unsigned_3 = '0;
  localparam bit unsigned [3:0] bit_unsigned_4 = '1;
  localparam bit unsigned [2:0][3:0] bit_unsigned_5 = '0;
  localparam bit unsigned [2:0][3:0] bit_unsigned_6 = '1;
  localparam bit unsigned [2:0][3:0] bit_unsigned_7 = '{1, 2, 3};
  localparam bit unsigned [2:0][3:0] bit_unsigned_8 = {4'd1, 4'd2, 4'd3};
  localparam bit signed [3:0] bit_signed_0 = 4'b0101;
  localparam bit signed [3:0] bit_signed_1 = 4'd5;
  localparam bit signed [3:0] bit_signed_2 = 5;
  localparam bit signed [3:0] bit_signed_3 = '0;
  localparam bit signed [3:0] bit_signed_4 = '1;
  localparam bit signed [2:0][3:0] bit_signed_5 = '0;
  localparam bit signed [2:0][3:0] bit_signed_6 = '1;
  localparam bit signed [2:0][3:0] bit_signed_7 = '{1, 2, 3};
  localparam bit signed [2:0][3:0] bit_signed_8 = {4'd1, 4'd2, 4'd3};

  localparam logic [3:0] logic_0 = 4'b0101;
  localparam logic [3:0] logic_1 = 4'd5;
  localparam logic [3:0] logic_2 = 5;
  localparam logic [3:0] logic_3 = '0;
  localparam logic [3:0] logic_4 = '1;
  localparam logic [2:0][3:0] logic_5 = '0;
  localparam logic [2:0][3:0] logic_6 = '1;
  localparam logic [2:0][3:0] logic_7 = '{1, 2, 3};
  localparam logic [2:0][3:0] logic_8 = {4'd1, 4'd2, 4'd3};
  localparam logic [2:0][3:0] logic_9 = 'X;
  localparam logic [2:0][3:0] logic_10 = 'Z;
  localparam logic unsigned [3:0] logic_unsigned_0 = 4'b0101;
  localparam logic unsigned [3:0] logic_unsigned_1 = 4'd5;
  localparam logic unsigned [3:0] logic_unsigned_2 = 5;
  localparam logic unsigned [3:0] logic_unsigned_3 = '0;
  localparam logic unsigned [3:0] logic_unsigned_4 = '1;
  localparam logic unsigned [2:0][3:0] logic_unsigned_5 = '0;
  localparam logic unsigned [2:0][3:0] logic_unsigned_6 = '1;
  localparam logic unsigned [2:0][3:0] logic_unsigned_7 = '{1, 2, 3};
  localparam logic unsigned [2:0][3:0] logic_unsigned_8 = {4'd1, 4'd2, 4'd3};
  localparam logic unsigned [2:0][3:0] logic_unsigned_9 = 'X;
  localparam logic unsigned [2:0][3:0] logic_unsigned_10 = 'Z;
  localparam logic signed [3:0] logic_signed_0 = 4'b0101;
  localparam logic signed [3:0] logic_signed_1 = 4'd5;
  localparam logic signed [3:0] logic_signed_2 = 5;
  localparam logic signed [3:0] logic_signed_3 = '0;
  localparam logic signed [3:0] logic_signed_4 = '1;
  localparam logic signed [2:0][3:0] logic_signed_5 = '0;
  localparam logic signed [2:0][3:0] logic_signed_6 = '1;
  localparam logic signed [2:0][3:0] logic_signed_7 = '{1, 2, 3};
  localparam logic signed [2:0][3:0] logic_signed_8 = {4'd1, 4'd2, 4'd3};
  localparam logic signed [2:0][3:0] logic_signed_9 = 'X;
  localparam logic signed [2:0][3:0] logic_signed_10 = 'Z;

  localparam reg [3:0] reg_0 = 4'b0101;
  localparam reg [3:0] reg_1 = 4'd5;
  localparam reg [3:0] reg_2 = 5;
  localparam reg [3:0] reg_3 = '0;
  localparam reg [3:0] reg_4 = '1;
  localparam reg [2:0][3:0] reg_9 = 'X;
  localparam reg [2:0][3:0] reg_10 = 'Z;
  localparam reg [2:0][3:0] reg_5 = '0;
  localparam reg [2:0][3:0] reg_6 = '1;
  localparam reg [2:0][3:0] reg_7 = '{1, 2, 3};
  localparam reg [2:0][3:0] reg_8 = {4'd1, 4'd2, 4'd3};
  localparam reg unsigned [3:0] reg_unsigned_0 = 4'b0101;
  localparam reg unsigned [3:0] reg_unsigned_1 = 4'd5;
  localparam reg unsigned [3:0] reg_unsigned_2 = 5;
  localparam reg unsigned [3:0] reg_unsigned_3 = '0;
  localparam reg unsigned [3:0] reg_unsigned_4 = '1;
  localparam reg unsigned [2:0][3:0] reg_unsigned_5 = '0;
  localparam reg unsigned [2:0][3:0] reg_unsigned_6 = '1;
  localparam reg unsigned [2:0][3:0] reg_unsigned_7 = '{1, 2, 3};
  localparam reg unsigned [2:0][3:0] reg_unsigned_8 = {4'd1, 4'd2, 4'd3};
  localparam reg unsigned [2:0][3:0] reg_unsigned_9 = 'X;
  localparam reg unsigned [2:0][3:0] reg_unsigned_10 = 'Z;
  localparam reg signed [3:0] reg_signed_0 = 4'b0101;
  localparam reg signed [3:0] reg_signed_1 = 4'd5;
  localparam reg signed [3:0] reg_signed_2 = 5;
  localparam reg signed [3:0] reg_signed_3 = '0;
  localparam reg signed [3:0] reg_signed_4 = '1;
  localparam reg signed [2:0][3:0] reg_signed_5 = '0;
  localparam reg signed [2:0][3:0] reg_signed_6 = '1;
  localparam reg signed [2:0][3:0] reg_signed_7 = '{1, 2, 3};
  localparam reg signed [2:0][3:0] reg_signed_8 = {4'd1, 4'd2, 4'd3};
  localparam reg signed [2:0][3:0] reg_signed_9 = 'X;
  localparam reg signed [2:0][3:0] reg_signed_10 = 'Z;
endpackage // }}} P_integralVectorPacked

package P_integralVectorUnpacked; // {{{
  localparam bit       bit_0  [1]   = '{1};
  localparam bit [2:0] bit_1  [1]   = '{3};
  localparam bit [2:0] bit_2  [0:0] = '{3};
  localparam bit       bit_3  [3]   = '{1, 1, 0};
  localparam bit       bit_4  [2:0] = '{1, 1, 0};
  localparam bit       bit_5  [0:2] = '{0, 1, 1};
  localparam bit [0:0] bit_6  [3]   = '{1, 1, 0};
  localparam bit [0:0] bit_7  [2:0] = '{1, 1, 0};
  localparam bit [0:0] bit_8  [0:2] = '{0, 1, 1};
  localparam bit [2:0] bit_9  [3]   = '{3, 2, 1};
  localparam bit [2:0] bit_10 [2:0] = '{3, 2, 1};
  localparam bit [2:0] bit_11 [0:2] = '{1, 2, 3};
  localparam bit unsigned       bit_unsigned_0  [1]   = '{1};
  localparam bit unsigned [2:0] bit_unsigned_1  [1]   = '{3};
  localparam bit unsigned [2:0] bit_unsigned_2  [0:0] = '{3};
  localparam bit unsigned       bit_unsigned_3  [3]   = '{1, 1, 0};
  localparam bit unsigned       bit_unsigned_4  [2:0] = '{1, 1, 0};
  localparam bit unsigned       bit_unsigned_5  [0:2] = '{0, 1, 1};
  localparam bit unsigned [0:0] bit_unsigned_6  [3]   = '{1, 1, 0};
  localparam bit unsigned [0:0] bit_unsigned_7  [2:0] = '{1, 1, 0};
  localparam bit unsigned [0:0] bit_unsigned_8  [0:2] = '{0, 1, 1};
  localparam bit unsigned [2:0] bit_unsigned_9  [3]   = '{3, 2, 1};
  localparam bit unsigned [2:0] bit_unsigned_10 [2:0] = '{3, 2, 1};
  localparam bit unsigned [2:0] bit_unsigned_11 [0:2] = '{1, 2, 3};
  localparam bit signed       bit_signed_0  [1]   = '{1};
  localparam bit signed [2:0] bit_signed_1  [1]   = '{3};
  localparam bit signed [2:0] bit_signed_2  [0:0] = '{3};
  localparam bit signed       bit_signed_3  [3]   = '{1, 1, 0};
  localparam bit signed       bit_signed_4  [2:0] = '{1, 1, 0};
  localparam bit signed       bit_signed_5  [0:2] = '{0, 1, 1};
  localparam bit signed [0:0] bit_signed_6  [3]   = '{1, 1, 0};
  localparam bit signed [0:0] bit_signed_7  [2:0] = '{1, 1, 0};
  localparam bit signed [0:0] bit_signed_8  [0:2] = '{0, 1, 1};
  localparam bit signed [2:0] bit_signed_9  [3]   = '{3, 2, 1};
  localparam bit signed [2:0] bit_signed_10 [2:0] = '{3, 2, 1};
  localparam bit signed [2:0] bit_signed_11 [0:2] = '{1, 2, 3};

  localparam logic       logic_0  [1]   = '{1};
  localparam logic [2:0] logic_1  [1]   = '{3};
  localparam logic [2:0] logic_2  [0:0] = '{3};
  localparam logic       logic_3  [3]   = '{1, 1, 0};
  localparam logic       logic_4  [2:0] = '{1, 1, 0};
  localparam logic       logic_5  [0:2] = '{0, 1, 1};
  localparam logic [0:0] logic_6  [3]   = '{1, 1, 0};
  localparam logic [0:0] logic_7  [2:0] = '{1, 1, 0};
  localparam logic [0:0] logic_8  [0:2] = '{0, 1, 1};
  localparam logic [2:0] logic_9  [3]   = '{3, 2, 1};
  localparam logic [2:0] logic_10 [2:0] = '{3, 2, 1};
  localparam logic [2:0] logic_11 [0:2] = '{1, 2, 3};
  localparam logic [2:0] logic_12 [3]   = '{'X, 'Z, 'X};
  localparam logic unsigned       logic_unsigned_0  [1]   = '{1};
  localparam logic unsigned [2:0] logic_unsigned_1  [1]   = '{3};
  localparam logic unsigned [2:0] logic_unsigned_2  [0:0] = '{3};
  localparam logic unsigned       logic_unsigned_3  [3]   = '{1, 1, 0};
  localparam logic unsigned       logic_unsigned_4  [2:0] = '{1, 1, 0};
  localparam logic unsigned       logic_unsigned_5  [0:2] = '{0, 1, 1};
  localparam logic unsigned [0:0] logic_unsigned_6  [3]   = '{1, 1, 0};
  localparam logic unsigned [0:0] logic_unsigned_7  [2:0] = '{1, 1, 0};
  localparam logic unsigned [0:0] logic_unsigned_8  [0:2] = '{0, 1, 1};
  localparam logic unsigned [2:0] logic_unsigned_9  [3]   = '{3, 2, 1};
  localparam logic unsigned [2:0] logic_unsigned_10 [2:0] = '{3, 2, 1};
  localparam logic unsigned [2:0] logic_unsigned_11 [0:2] = '{1, 2, 3};
  localparam logic unsigned [2:0] logic_unsigned_12 [3]   = '{'X, 'Z, 'Z};
  localparam logic signed       logic_signed_0  [1]   = '{1};
  localparam logic signed [2:0] logic_signed_1  [1]   = '{3};
  localparam logic signed [2:0] logic_signed_2  [0:0] = '{3};
  localparam logic signed       logic_signed_3  [3]   = '{1, 1, 0};
  localparam logic signed       logic_signed_4  [2:0] = '{1, 1, 0};
  localparam logic signed       logic_signed_5  [0:2] = '{0, 1, 1};
  localparam logic signed [0:0] logic_signed_6  [3]   = '{1, 1, 0};
  localparam logic signed [0:0] logic_signed_7  [2:0] = '{1, 1, 0};
  localparam logic signed [0:0] logic_signed_8  [0:2] = '{0, 1, 1};
  localparam logic signed [2:0] logic_signed_9  [3]   = '{3, 2, 1};
  localparam logic signed [2:0] logic_signed_10 [2:0] = '{3, 2, 1};
  localparam logic signed [2:0] logic_signed_11 [0:2] = '{1, 2, 3};
  localparam logic signed [2:0] logic_signed_12 [3]   = '{'X, 'Z, 'Z};

  localparam reg       reg_0  [1]   = '{1};
  localparam reg [2:0] reg_1  [1]   = '{3};
  localparam reg [2:0] reg_2  [0:0] = '{3};
  localparam reg       reg_3  [3]   = '{1, 1, 0};
  localparam reg       reg_4  [2:0] = '{1, 1, 0};
  localparam reg       reg_5  [0:2] = '{0, 1, 1};
  localparam reg [0:0] reg_6  [3]   = '{1, 1, 0};
  localparam reg [0:0] reg_7  [2:0] = '{1, 1, 0};
  localparam reg [0:0] reg_8  [0:2] = '{0, 1, 1};
  localparam reg [2:0] reg_9  [3]   = '{3, 2, 1};
  localparam reg [2:0] reg_10 [2:0] = '{3, 2, 1};
  localparam reg [2:0] reg_11 [0:2] = '{1, 2, 3};
  localparam reg [2:0] reg_12 [3]   = '{'X, 'Z, 'X};
  localparam reg unsigned       reg_unsigned_0  [1]   = '{1};
  localparam reg unsigned [2:0] reg_unsigned_1  [1]   = '{3};
  localparam reg unsigned [2:0] reg_unsigned_2  [0:0] = '{3};
  localparam reg unsigned       reg_unsigned_3  [3]   = '{1, 1, 0};
  localparam reg unsigned       reg_unsigned_4  [2:0] = '{1, 1, 0};
  localparam reg unsigned       reg_unsigned_5  [0:2] = '{0, 1, 1};
  localparam reg unsigned [0:0] reg_unsigned_6  [3]   = '{1, 1, 0};
  localparam reg unsigned [0:0] reg_unsigned_7  [2:0] = '{1, 1, 0};
  localparam reg unsigned [0:0] reg_unsigned_8  [0:2] = '{0, 1, 1};
  localparam reg unsigned [2:0] reg_unsigned_9  [3]   = '{3, 2, 1};
  localparam reg unsigned [2:0] reg_unsigned_10 [2:0] = '{3, 2, 1};
  localparam reg unsigned [2:0] reg_unsigned_11 [0:2] = '{1, 2, 3};
  localparam reg unsigned [2:0] reg_unsigned_12 [3]   = '{'X, 'Z, 'Z};
  localparam reg signed       reg_signed_0  [1]   = '{1};
  localparam reg signed [2:0] reg_signed_1  [1]   = '{3};
  localparam reg signed [2:0] reg_signed_2  [0:0] = '{3};
  localparam reg signed       reg_signed_3  [3]   = '{1, 1, 0};
  localparam reg signed       reg_signed_4  [2:0] = '{1, 1, 0};
  localparam reg signed       reg_signed_5  [0:2] = '{0, 1, 1};
  localparam reg signed [0:0] reg_signed_6  [3]   = '{1, 1, 0};
  localparam reg signed [0:0] reg_signed_7  [2:0] = '{1, 1, 0};
  localparam reg signed [0:0] reg_signed_8  [0:2] = '{0, 1, 1};
  localparam reg signed [2:0] reg_signed_9  [3]   = '{3, 2, 1};
  localparam reg signed [2:0] reg_signed_10 [2:0] = '{3, 2, 1};
  localparam reg signed [2:0] reg_signed_11 [0:2] = '{1, 2, 3};
  localparam reg signed [2:0] reg_signed_12 [3]   = '{'X, 'Z, 'Z};
endpackage // }}} P_integralVectorUnpacked
