module TestModule
( output my_enum_t d
, output var my_struct_t e, f
);
endmodule