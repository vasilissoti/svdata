module mh9(output signed [5:0] x);
endmodule