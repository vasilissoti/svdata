module mh1 (integer x); 
endmodule