module TestModule
( a, [FOO-1:0] b
, wire [FOO-1:0] c [FOO] [FOO-1:0], int d
, logic e [FOO-1:0], f
, string g
, inout unsigned h
, inout tri integer unsigned i
);
endmodule