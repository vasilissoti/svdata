module mh3 ([5:0] x);
endmodule