module mh7 (output x);
endmodule