module TestModule
( input var signed [FOO-1:0] a [FOO] [FOO-1:0], b
, input var signed c, var reg signed d
, input var logic signed e [FOO-1:0]
, input var integer signed f
);
endmodule