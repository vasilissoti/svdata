module TestModule
( output signed [FOO-1:0] a [FOO] [FOO-1:0], b
, output wire logic signed [FOO-1:0] c, wire reg signed d
, output tri integer signed e
);
endmodule