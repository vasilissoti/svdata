module mh17(output var x, input y);
endmodule