module TestModule
( signed a, signed [FOO-1:0] b
, wire signed [FOO-1:0] c, int signed d
, logic signed e [DOO-1:0], f
, inout signed g
, inout tri integer signed h
);
endmodule