module mh16(input var integer x, wire y);
endmodule