module TestModule
#(parameter a = 8'sb10101010 + 6'sb10101010,
  parameter b = 4'b1000 + 3.5 -2,
  parameter c = -2 + 3 + 5 + 8'sb10101010,
  parameter e = -2 + 3 + 5 + 8'b10101010,
  parameter f = -2.5 + 3.5 + 4.5)
(); 
endmodule