module mh12(ref x [5:0]);
endmodule