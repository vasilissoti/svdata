module TestModule
( input var [FOO-1:0] a [FOO] [FOO-1:0], b
, input var c, var reg d
, input var logic e [FOO-1:0]
, input var string f
, input var integer unsigned g
);
endmodule