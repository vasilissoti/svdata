module TestModule
( inout my_enum_t d
, inout wire my_struct_t e, f
);
endmodule