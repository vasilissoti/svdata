module TestModule
#(localparam a = 8'sb10101010, 
  localparam logic signed [3:0] b = 4'b1000,
  localparam c = 7.5, d = 5,
  localparam e = "hello")
(); 
endmodule