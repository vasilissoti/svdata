module TestModule
#(localparam a = (8'sb10101010 + "hello") /* A0 */, b = 3, // A1
parameter /* B0 */ c = 1 /* B1 */, d = 6, e)
(); 
endmodule