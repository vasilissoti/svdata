module mh2 (inout integer x);
endmodule