module TestModule
  #(/*pre*/ a /*post*/
  , /*pre*/ b /*id/eq*/ = /*eq/val*/ 5 /*post*/
  , /*pre*/ int /*ty/id*/ c /*post*/
  , /*pre*/ int /*ty/id*/ d /* id/eq */ = /*eq/val*/ 5 /*post*/)
  ();
endmodule