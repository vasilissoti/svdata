module TestModule
( input signed [FOO-1:0] a, b
, input wire signed [FOO-1:0] c, reg signed d
, input logic signed e [FOO-1:0]
, input tri integer signed f
);
endmodule