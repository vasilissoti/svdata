module Loo
( a, signed b
);
endmodule