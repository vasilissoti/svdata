package TestPackage;
  parameter a = 8'sb10101010;
  parameter logic signed [3:0] b = 4'b1000;
  parameter e = 7.5, f = 5;
  parameter g = "hello";
endpackage