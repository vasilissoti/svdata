package TestPackage;
  localparam a = 8'sb10101010;
  localparam logic signed [3:0] b = 4'b1000;
  localparam e = 7.5, f = 5;
  localparam g = "hello";
endpackage