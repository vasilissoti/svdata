package foo;
endpackage

module Foo();
endmodule

package bar;
endpackage

module Bar();
endmodule
