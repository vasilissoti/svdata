module TestModule
#(integer a = 8'sb10101010, 
  logic signed [3:0] b = 4'b1000, c [4:0],
  real e = 7.5, 
  integer f = 5,
  string g = "hello")
(); 
endmodule